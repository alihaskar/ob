//========================================================================== //
// Copyright (c) 2020, Stephen Henry
// All rights reserved.
//
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// * Redistributions of source code must retain the above copyright notice, this
//   list of conditions and the following disclaimer.
//
// * Redistributions in binary form must reproduce the above copyright notice,
//   this list of conditions and the following disclaimer in the documentation
//   and/or other materials provided with the distribution.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
// ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
// INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
// CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.
//========================================================================== //

`include "ob_pkg.vh"
`include "ob_cntrl_pkg.vh"

module ob_cntrl_dec (
  // ======================================================================== //
  // Encoded instruction:
    input ob_cntrl_pkg::inst_t                    inst

  // ======================================================================== //
  // Decoded micro-code:
  , output ob_cntrl_pkg::ucode_t                  ucode
);

  function automatic ob_cntrl_pkg::ucode_t decode__nop(); begin
    return '0;
  end endfunction


  function automatic ob_cntrl_pkg::ucode_t decode__search_result_common(
    ob_pkg::search_result_t sr); begin
    ob_pkg::result_trade_t trade;
    ob_cntrl_pkg::ucode_t uc;

    // Microcode defaults:
    uc                  = '0;

    // Emit output response
    uc.rsp_vld          = 'b1;

    uc.rsp              = '0;
    // Trade has no originator command therefore UID is set as '1 to indicate
    // that this response was internally generated by the matching engine.
    uc.rsp.uid          = '1;
    uc.rsp.status       = ob_pkg::S_Okay;

    // Form trade response oprand.
    trade               = '0;
    trade.bid_uid       = sr.bid_uid;
    trade.ask_uid       = sr.ask_uid;
    trade.quantity      = sr.quantity;

    uc.rsp.result.trade = trade;

    return uc;
  end endfunction


  function automatic ob_cntrl_pkg::ucode_t decode__lm_ask_lm_bid(
    ob_pkg::search_result_t sr); begin
    ob_cntrl_pkg::ucode_t uc = decode__search_result_common(sr);

    case ({sr.bid_consumed, sr.ask_consumed}) inside
      2'b10: begin
        // Limit bid head has been consumed by current match
        uc.lm_bid_pop             = 'b1;
        // Limit ask head update.
        uc.lm_ask_update_vld      = 'b1;
        uc.lm_ask_update          = '0;
        uc.lm_ask_update.uid      = sr.ask_uid;
        uc.lm_ask_update.price    = sr.ask_price;
        uc.lm_ask_update.quantity = sr.remainder;
      end
      2'b01: begin
        // Limit ask head has been consumed by current match
        uc.lm_ask_pop = 'b1;
        // Limit bid head update.
        uc.lm_bid_update_vld      = 'b1;
        uc.lm_bid_update          = '0;
        uc.lm_bid_update.uid      = sr.bid_uid;
        uc.lm_bid_update.price    = sr.bid_price;
        uc.lm_bid_update.quantity = sr.remainder;
      end
      2'b11: begin
        // Both bid/ask heads have been consumed by current match.
        uc.lm_bid_pop = 'b1;
        uc.lm_ask_pop = 'b1;
      end
      default: begin
        // Otherwise,
      end
    endcase
    return uc;
  end endfunction


  function automatic ob_cntrl_pkg::ucode_t decode__lm_ask_mk_bid(
    ob_pkg::search_result_t sr); begin
    ob_cntrl_pkg::ucode_t uc = decode__search_result_common(sr);
    return uc;
  end endfunction

  function automatic ob_cntrl_pkg::ucode_t decode__mk_ask_lm_bid(
    ob_pkg::search_result_t sr); begin
    ob_cntrl_pkg::ucode_t uc = decode__search_result_common(sr);
    return uc;
  end endfunction

  function automatic ob_cntrl_pkg::ucode_t decode__mk_ask_mk_bid(
    ob_pkg::search_result_t sr); begin
    ob_cntrl_pkg::ucode_t uc = decode__search_result_common(sr);
    return uc;
  end endfunction

  function automatic ob_cntrl_pkg::ucode_t decode__emit_rsp(
    ob_pkg::uid_t uid, ob_pkg::status_t status); begin

    ob_cntrl_pkg::ucode_t uc = '0;
    // Issue response:
    uc.rsp_vld               = 'b1;
    // Form response packet:
    uc.rsp                   = '0;
    uc.rsp.uid               = uid;
    uc.rsp.status            = status;
    uc.rsp.result            = '0;
    return uc;
  end endfunction

  function automatic ob_cntrl_pkg::ucode_t decode__push_table(
    ob_pkg::cmd_t cmd, ob_cntrl_pkg::table_id_t id); begin
    ob_cntrl_pkg::ucode_t uc;

    uc = '0;

    // Issue table command
    case (id)
      ob_cntrl_pkg::TBL_ID__LM_ASK: begin
        // Issue insert command:
        uc.lm_ask_insert              = 'b1;
        // Form insert payload:
        uc.lm_ask_insert_tbl          = '0;
        uc.lm_ask_insert_tbl.uid      = cmd.uid;
        uc.lm_ask_insert_tbl.quantity = cmd.quantity;
        uc.lm_ask_insert_tbl.price    = cmd.price;
      end
      ob_cntrl_pkg::TBL_ID__LM_BID: begin
        // Issue insert command:
        uc.lm_bid_insert              = 'b1;
        // Form insert payload:
        uc.lm_bid_insert_tbl          = '0;
        uc.lm_bid_insert_tbl.uid      = cmd.uid;
        uc.lm_bid_insert_tbl.quantity = cmd.quantity;
        uc.lm_bid_insert_tbl.price    = cmd.price;
      end
      ob_cntrl_pkg::TBL_ID__MK_ASK: begin
        // Issue insert command:
        uc.mk_ask_insert              = 'b1;
        // Form insert payload:
        uc.mk_ask_insert_tbl          = '0;
        uc.mk_ask_insert_tbl.uid      = cmd.uid;
        uc.mk_ask_insert_tbl.quantity = cmd.quantity;
        uc.mk_ask_insert_tbl.price    = cmd.price;
      end
      ob_cntrl_pkg::TBL_ID__MK_BID: begin
        // Issue insert command:
        uc.mk_bid_insert              = 'b1;
        // Form insert payload:
        uc.mk_bid_insert_tbl          = '0;
        uc.mk_bid_insert_tbl.uid      = cmd.uid;
        uc.mk_bid_insert_tbl.quantity = cmd.quantity;
        uc.mk_bid_insert_tbl.price    = cmd.price;
      end
      default: begin
        // Invalid table destination.
      end
    endcase // case (id)

    // Issue response
    uc.rsp_vld    = 'b1;

    // Response message:
    uc.rsp        = '0;
    uc.rsp.uid    = cmd.uid;
    uc.rsp.status = ob_pkg::S_Okay;

    return uc;
  end endfunction

  function automatic ob_cntrl_pkg::ucode_t decode__pop_table(
    ob_cntrl_pkg::table_id_t id); begin

    ob_cntrl_pkg::ucode_t uc;

    uc = '0;

    // Issue table command
    case (id)
      ob_cntrl_pkg::TBL_ID__LM_ASK: begin
      end
      ob_cntrl_pkg::TBL_ID__LM_BID: begin
      end
      ob_cntrl_pkg::TBL_ID__MK_ASK: begin
      end
      ob_cntrl_pkg::TBL_ID__MK_BID: begin
      end
      default: begin
        // Invalid table destination.
      end
    endcase // case (id)

    // Issue response
    uc.rsp_vld = 'b1;


    return uc;
  end endfunction

  // ------------------------------------------------------------------------ //
  //
  always_comb begin : decode_PROC

    ucode = decode__nop();

    case (inst.opcode)
      ob_cntrl_pkg::OP_NOP: begin
      end
      ob_cntrl_pkg::OP_SEARCH_RESULT: begin
        ob_pkg::search_result_t sr = inst.oprand.search_result.sr;

        case ({// Limit Ask <-> Limit Bid
               sr.lm_ask_lm_bid,
               // Limit Ask <-> Market Bid
               sr.lm_ask_mk_bid,
               // Market Ask <-> Limit Bid
               sr.mk_ask_lm_bid,
               // Market Ask <-> Market Bid
               sr.mk_ask_mk_bid}) inside
          4'b1???: begin
            // Trade on Limit Ask (Sell) <-> Limit Bid (Buy)
            ucode = decode__lm_ask_lm_bid(sr);
          end
          4'b01??: begin
            // Trade on Limit Ask (Sell) <-> Market Bid (Buy)
            ucode = decode__lm_ask_mk_bid(sr);
          end
          4'b001?: begin
            // Trade on Market Ask (Sell) <-> Limit Bid (Buy)
            ucode = decode__mk_ask_lm_bid(sr);
          end
          4'b0001: begin
            // Trade on Market Ask (Sell) <-> Market Bid (Buy)
            ucode = decode__mk_ask_mk_bid(sr);
          end
          default: begin
            // Error, a match should have been detected.
            ucode = decode__nop();
          end
        endcase // case ({...

      end // case: ob_cntrl_pkg::OP_SEARCH_RESULT
      ob_cntrl_pkg::OP_EMIT_RSP: begin
        // Issue response notification:
        ucode = decode__emit_rsp(
          .uid(inst.oprand.emit_rsp.uid), .status(inst.oprand.emit_rsp.status));
      end
      ob_cntrl_pkg::OP_PUSH_TABLE: begin
        ucode = decode__push_table(
          .cmd(inst.oprand.push_table.cmd), .id(inst.oprand.push_table.table_id));
      end
      ob_cntrl_pkg::OP_POP_TABLE: begin
        ucode = decode__pop_table(.id(inst.oprand.pop_table.table_id));
      end
      default: begin
        // Unknown opcode (raise error condition?).
      end
    endcase // case (inst.opcode)

  end

endmodule // ob_cntrl_dec
